// Simple example: variable initialization and finish
module Top;
  int x = 42;
  initial $finish;
endmodule
