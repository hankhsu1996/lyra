module Test;
  int a, b, c;
  initial begin
    a = 1;
    b = 2;
    c = a + b;
  end
endmodule
